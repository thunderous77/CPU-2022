`include "D:/Sam/program/CPU-2022/riscv/src/defines.v"

module ROB(
    input wire clk,
    input wire rst,
    input wire rdy,

    // 
);

endmodule